package apb_test_pkg;

    import uvm_pkg::*;   //import the uvm package library

    import apb_bridge_agent_pkg::*;  //import the apb bridge/master agent package
    
    import apb_slave_agent_pkg::*;   //import the apb slave agent package
    
    import apb_environment_pkg::*;           //import the apb environment package
    
    `include "uvm_macros.svh"   //include the uvm macros file
    
    `include "apb_config.svh"   //include apb configuration file

    `include "apb_slave_seqc.svh"
    `include "apb_bridge_seqc.svh"
    `include "apb_virtual_seqc.svh"
    `include "apb_virtual_seqc_write.svh"

    `include "apb_test_base.svh"  //include apb_test_base file
    `include "apb_test_write.svh"
    
endpackage:apb_test_pkg
