package apb_slave_agent_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"
    `include "apb_config.svh"   //include apb configuration file
    `include "apb_slave_config_obj.svh"
    `include "apb_slave_seq_item.svh"
    `include "apb_storage_component.svh"
    `include "apb_slave_sequencer.svh"
    `include "apb_slave_drv.svh"
    `include "apb_slave_agent.svh"

endpackage
