`define ADDR_BUS_WIDTH 32

`define DATA_BUS_BYTES 4

`define NO_OF_SLAVE_ON_BUS 1
