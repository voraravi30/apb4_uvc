package apb_environment_pkg;

    import uvm_pkg::*;
    import apb_bridge_agent_pkg::*;
    import apb_slave_agent_pkg::*;

    `include "uvm_macros.svh"
    `include "apb_config.svh"   //include apb configuration file

    `include "apb_env_config.svh"
    `include "apb_predictor.svh"
    `include "apb_comparator.svh"
    `include "apb_scoreboard.svh"
    `include "apb_bus_monitor.svh"
    `include "apb_coverage.svh"
    `include "apb_virtual_sequencer.svh"
    `include "apb_environment.svh"

endpackage
