package apb_sequence_pkg;

    import uvm_pkg::*;
    import apb_bridge_agent_pkg::*;
    import apb_slave_agent_pkg::*;

    `include "uvm_macros.svh"
    `include "apb_config.svh"   //include apb configuration file
    `include "apb_slave_sequence.svh"
    `include "apb_bridge_sequence.svh"
    `include "apb_virtual_sequence.svh"

endpackage:apb_sequence_pkg
